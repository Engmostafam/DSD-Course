/*
*/ 

module stpmtr (/*AUTOARG*/);

   
 
endmodule // stpmtr


