module pnser (/*AUTOARG*/);
 
endmodule // pnser

